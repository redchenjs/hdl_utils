/*
 * ahb2mmio.sv
 *
 *  Created on: 2023-08-09 22:26
 *      Author: Jack Chen <redchenjs@live.com>
 */

`timescale 1 ns / 1 ps

import ahb_enum::*;

module ahb2mmio #(
    parameter A_WIDTH = 32,
    parameter D_WIDTH = 32
) (
    input logic hclk_i,
    input logic hresetn_i,

    // ahb port
    input logic               hsel_i,
    input logic [A_WIDTH-1:0] haddr_i,
    input logic         [3:0] hprot_i,
    input logic         [2:0] hsize_i,
    input logic         [1:0] htrans_i,
    input logic         [2:0] hburst_i,
    input logic               hwrite_i,
    input logic [D_WIDTH-1:0] hwdata_i,

    output logic         [1:0] hresp_o,
    output logic               hready_o,
    output logic [D_WIDTH-1:0] hrdata_o,

    // mmio port
    output logic [D_WIDTH/8-1:0] wr_en_o,
    output logic   [A_WIDTH-1:0] wr_addr_o,
    output logic   [D_WIDTH-1:0] wr_data_o,

    output logic               rd_en_o,
    output logic [A_WIDTH-1:0] rd_addr_o,
    input  logic [D_WIDTH-1:0] rd_data_i
);

logic                 hsel_r;
logic [D_WIDTH/8-1:0] hsel_w;
logic   [A_WIDTH-1:0] haddr_w;

logic [D_WIDTH/8-1:0] [$clog2(D_WIDTH/8):0] [D_WIDTH/8-1:0] hsel_mux;

assign wr_en_o   = hsel_w;
assign wr_addr_o = haddr_w;
assign wr_data_o = hwdata_i;

assign rd_en_o   = hsel_r;
assign rd_addr_o = haddr_i;

assign hresp_o  = AHB_RESP_OKAY;
assign hready_o = 'b1;
assign hrdata_o = rd_data_i;

generate
    genvar i;

    for (i = 0; i < $clog2(D_WIDTH/8)+1; i++) begin: gen_en_sel
        genvar j;

        for (j = 0; j < D_WIDTH/8; j++) begin: gen_en_bit
            genvar k;

            for (k = 0; k < D_WIDTH/8; k++) begin: gen_en_sft
                assign hsel_mux[k][i][j] =(j < ((1 << i) + k)) & (j >= k);
            end
        end
    end
endgenerate

always_comb begin
    case (htrans_i)
        AHB_TRANS_IDLE,
        AHB_TRANS_BUSY: begin
            hsel_r = 'b0;
        end
        AHB_TRANS_NONSEQ,
        AHB_TRANS_SEQ: begin
            hsel_r = hsel_i & !hwrite_i;
        end
        default: begin
            hsel_r = 'b0;
        end
    endcase
end

always_ff @(posedge hclk_i or negedge hresetn_i)
begin
    if (!hresetn_i) begin
        hsel_w  <= 'b0;
        haddr_w <= 'b0;
    end else begin
        case (htrans_i)
            AHB_TRANS_IDLE,
            AHB_TRANS_BUSY: begin
                hsel_w  <= 'b0;
                haddr_w <= 'b0;
            end
            AHB_TRANS_NONSEQ,
            AHB_TRANS_SEQ: begin
                hsel_w  <= hsel_i & hwrite_i ? hsel_mux[haddr_i[$clog2(D_WIDTH/8)-1:0]][hsize_i] : 'b0;
                haddr_w <= haddr_i;
            end
            default: begin
                hsel_w  <= 'b0;
                haddr_w <= 'b0;
            end
        endcase
    end
end

endmodule
